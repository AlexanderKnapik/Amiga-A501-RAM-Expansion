module a501(
	    input [8:0] addressIn,
	    input [3:0] rtcAddress,
	    inout [3:0] rtcData,
	    output [17:0] addressOut
)

 
      
      
endmodule // a501

